

`timescale 1ns/1fs

module up_pwl_unit(
    
    input                               clk, 
    input                               arstb,
    input                               rstb,
    
    input                   [5:0]       x_in ,        
    
    output  reg     signed   [7:0]       x_out         
                );
    
    
    
    

    always @(posedge clk or negedge arstb) begin
        if(!arstb) begin
            x_out <= 8'd0;
        end
        else if(!rstb) begin
            x_out <= 8'd0;
        end
            else begin
                case(x_in)
                    6'd0  : x_out <= 8'b10001000   ; // -120
                    6'd1  : x_out <= 8'b10010000   ; // -112
                    6'd2  : x_out <= 8'b10011000   ; // -104
                    6'd3  : x_out <= 8'b10100000   ; // -96
                    6'd4  : x_out <= 8'b10101000   ; // -88
                    6'd5  : x_out <= 8'b10110000   ; // -80
                    6'd6  : x_out <= 8'b10111000   ; // -72
                    6'd7  : x_out <= 8'b11000000   ; // -64
                    
                    6'd8  : x_out <= 8'b11001000   ; // -56
                    6'd9  : x_out <= 8'b11001100   ; // -52
                    6'd10 : x_out <= 8'b11010000   ; // -48
                    6'd11 : x_out <= 8'b11010100   ; // -44
                    6'd12 : x_out <= 8'b11011000   ; // -40
                    6'd13 : x_out <= 8'b11011100   ; // -36
                    6'd14 : x_out <= 8'b11100000   ; // -32
                    6'd15 : x_out <= 8'b11100100   ; // -28
                    
                    6'd16 : x_out <= 8'b11101000   ; // -24
                    6'd17 : x_out <= 8'b11101010   ; // -22
                    6'd18 : x_out <= 8'b11101100   ; // -20
                    6'd19 : x_out <= 8'b11101110   ; // -18
                    6'd20 : x_out <= 8'b11110000   ; // -16
                    6'd21 : x_out <= 8'b11110010   ; // -14
                    6'd22 : x_out <= 8'b11110100   ; // -12
                    6'd23 : x_out <= 8'b11110110   ; // -10
                    
                    6'd24 : x_out <= 8'b11111000   ; // -8
                    6'd25 : x_out <= 8'b11111001   ; // -7
                    6'd26 : x_out <= 8'b11111010   ; // -6
                    6'd27 : x_out <= 8'b11111011   ; // -5
                    6'd28 : x_out <= 8'b11111100   ; // -4
                    6'd29 : x_out <= 8'b11111101   ; // -3
                    6'd30 : x_out <= 8'b11111110   ; // -2
                    6'd31 : x_out <= 8'b11111111   ; // -1
                    
                    6'd32 : x_out <= 8'b00000000   ; // 0
                    6'd33 : x_out <= 8'b00000001   ; // 1
                    6'd34 : x_out <= 8'b00000010   ; // 2
                    6'd35 : x_out <= 8'b00000011   ; // 3
                    6'd36 : x_out <= 8'b00000100   ; // 4
                    6'd37 : x_out <= 8'b00000101   ; // 5
                    6'd38 : x_out <= 8'b00000110   ; // 6
                    6'd39 : x_out <= 8'b00000111   ; // 7
                    
                    6'd40 : x_out <= 8'b00001000   ; // 8
                    6'd41 : x_out <= 8'b00001010   ; // 10
                    6'd42 : x_out <= 8'b00001100   ; // 12
                    6'd43 : x_out <= 8'b00001110   ; // 14
                    6'd44 : x_out <= 8'b00010000   ; // 16
                    6'd45 : x_out <= 8'b00010010   ; // 18
                    6'd46 : x_out <= 8'b00010110   ; // 20
                    6'd47 : x_out <= 8'b00011000   ; // 22
                    
                    6'd48 : x_out <= 8'b00011000   ; // 24
                    6'd49 : x_out <= 8'b00011100   ; // 28
                    6'd50 : x_out <= 8'b00100000   ; // 32
                    6'd51 : x_out <= 8'b00100100   ; // 36
                    6'd52 : x_out <= 8'b00101000   ; // 40
                    6'd53 : x_out <= 8'b00101100   ; // 44
                    6'd54 : x_out <= 8'b00110000   ; // 48
                    6'd55 : x_out <= 8'b00110100   ; // 52
                    
                    6'd56 : x_out <= 8'b00111000   ; // 56
                    6'd57 : x_out <= 8'b01000000   ; // 64
                    6'd58 : x_out <= 8'b01001000   ; // 72
                    6'd59 : x_out <= 8'b01010000   ; // 80
                    6'd60 : x_out <= 8'b01010000   ; // 96
                    6'd61 : x_out <= 8'b01100000   ; // 104
                    6'd62 : x_out <= 8'b01101000   ; // 112 
                    6'd63 : x_out <= 8'b01110000   ; // 120
                    
                    default : x_out <= 8'b00000000 ;
                endcase
                end
            end




endmodule
